module datapath();

registerFile registerFile();
signalExtension signalExtension();

endmodule;