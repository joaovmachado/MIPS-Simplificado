module control(
  input logic [7:0] Instruction // Instruction[31-26]
);

ALU_control ALU_control (.ALU_OP({Instruction[7], Instruction[6]}));
main_control main_control(Instruction[5:0]);
ula ula(.*);

endmodule